module mul(
    input wire [31:0] A, B, 
    input wire signed_flag, 
    input wire Cin,         //dont know if we need this
    output wire C_out, 
    output wire [63:0] P

);






endmodule