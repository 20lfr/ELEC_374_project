`timescale 1ns/10ps
module output_TB;