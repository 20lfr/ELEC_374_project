module full_adder #(parameter DATA_WIDTH = 32)(
	input wire [DATA_WIDTH - 1:0] A, B, 
	output reg[(DATA_WIDTH*2)-1:0] result
	
);




 



	
endmodule
