module CON_FF (
    input wire IR[31:0], BusMuxOut[31:0]; //data in from IR and Bus
    output wire toControl[31:0];          //output to control signals, must also include interaction
);                                        //with PC.+



    
endmodule