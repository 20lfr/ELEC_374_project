module Control(
    
);


endmodule