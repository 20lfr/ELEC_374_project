module CLA_add #(parameter DATA_WIDTH = 32)(
	input reg [DATA_WIDTH - 1:0] A, B, 
	output reg[(DATA_WIDTH*2)-1:0] result
	
);






	
endmodule
