module decoder4to16(
    input wire [3:0] in,  // 4-bit input
    output wire [15:0] out // 16-bit output
);

assign out = (in == 4'b0000) ? 16'b0000_0000_0000_0001 :
             (in == 4'b0001) ? 16'b0000_0000_0000_0010 :
             (in == 4'b0010) ? 16'b0000_0000_0000_0100 :
             (in == 4'b0011) ? 16'b0000_0000_0000_1000 :
             (in == 4'b0100) ? 16'b0000_0000_0001_0000 :
             (in == 4'b0101) ? 16'b0000_0000_0010_0000 :
             (in == 4'b0110) ? 16'b0000_0000_0100_0000 :
             (in == 4'b0111) ? 16'b0000_0000_1000_0000 :
             (in == 4'b1000) ? 16'b0000_0001_0000_0000 :
             (in == 4'b1001) ? 16'b0000_0010_0000_0000 :
             (in == 4'b1010) ? 16'b0000_0100_0000_0000 :
             (in == 4'b1011) ? 16'b0000_1000_0000_0000 :
             (in == 4'b1100) ? 16'b0001_0000_0000_0000 :
             (in == 4'b1101) ? 16'b0010_0000_0000_0000 :
             (in == 4'b1110) ? 16'b0100_0000_0000_0000 :
                               16'b1000_0000_0000_0000;

endmodule
